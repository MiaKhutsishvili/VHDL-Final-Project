----------------------------------------------------------------------------------
-- Kimia Khoodsiyani & Maral Torabi
-- 40223030            40223019

-- Create Date:    14:11:14 08/05/2025 
-- Module Name:    ALU - Behavioral 
-- Project Name: 	 Logical Circuits Final Project
-- Description:    This module is a simple calculator
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.Packages.All;

entity ALU is
    Port ( InPack : in  data_packet;
			  PackMode : in  packet_type;	
			  
			  SendToRam : out data_packet;
			  ReadResponse : in data_packet;
			  Finish : inout STD_LOGIC; 			-- Is 1 when the process is done.
			  
			  Enable : in STD_LOGIC;				-- Alu is On only when we are in Alu Mode.
			  Error : out STD_LOGIC;
			  RST : in STD_LOGIC;
			  clk : in STD_LOGIC
			 );
end ALU;

architecture Behavioral of ALU is	
	
	function Operator(In1, In2: signed(7 downto 0); operate : Alu_Operation) return byte is
	begin
		case operate is
			when Add => 
				return std_logic_vector(In1 + In2);
			when Sub => 
				return std_logic_vector(In1 - In2);
			when BitwiseOr => 
				return std_logic_vector(In1 or In2);		-- Bitwise or for signed = direct or
			when BitwiseAnd => 
				return std_logic_vector(In1 and In2);		-- Bitwise and for signed = direct and
			when others =>
				return "00000000";
		end case;
	end function;
	
	signal operation : Alu_Operation;
	---
	signal DataI : byte := (others => '0');
	signal DataII : byte := (others => '0');
		
	signal DestinationAddress : byte;
	signal ArrayLength : integer range 0 to 32 := 0;
	signal ArrayIndPusher : integer range 0 to 31 := 0;
	
	signal ReadArray : alu_read_cash_array := (others => (others => '0'));
		
	signal Step : integer := 0;
	
begin
	
	process(clk)
		-- Ram Interaction
		variable mode : byte := (others => '0');
		variable RamAddress : byte := (others => '0');								-- The Address given to the ram
		variable RamDataToWrite : byte := (others => '0');
		variable AddressI : byte := (others => '0');
		variable AddressII : byte := (others => '0');
		variable AddAddressII : byte := (others => '0');
		
		-- Calculator Interaction		
		
	begin
		if rising_edge(clk) then
			Error <= '0';
			if RST = '1' then
				Error <= '0';
				Step <= 0;
				DataI <= (others => '0');
				DataII <= (others => '0');
				DestinationAddress <= (others => '0');
				ArrayLength <= 0;
				ArrayIndPusher <= 0;
				ReadArray <= (others => (others => '0'));
				Finish <= '1';
			elsif Enable = '1' then
				if (Finish = '1') then				-- 1 * Clk -> 
					Finish <= '0';		
					case InPack(0)(1 downto 0) is 
						when "00" =>
							operation <= Add;
						when "01" => 
							operation <= Sub;
						when "10" => 
							operation <= BitwiseOr;
						when "11" =>
							operation <= BitwiseAnd;
						when others =>
					end case;			
				end if;
				
				case PackMode is 
					when Operand_Alu => -- 3 Clocks
						if Step = 0 then							-- Clock 0 till 1
							DestinationAddress <= InPack(3);
							AddressI := InPack(1);
							RamAddress := AddressI;
							mode := "00001111";
						elsif Step = 1 then						-- Clock 1 till 2
							DataI <= ReadResponse(1);
							AddressII := InPack(2);
							RamAddress := AddressII;
							mode := "00001111";
						elsif Step = 2 then						-- Clock 2 till 3
							--DataII <= ReadResponse(1);
							RamDataToWrite := Operator(signed(DataI), signed(ReadResponse(1)), Operation);
							RamAddress := DestinationAddress;
							mode := "11110000";
							Step <= -1;							-- Will + 1
							Finish <= '1';
						end if;
							
					when Immediate_Alu =>
						if Step = 0 then							-- Clock 0 till 1
							DataII <= InPack(2);
							DestinationAddress <= InPack(3);
							AddressI := InPack(1);
							RamAddress := AddressI;
							mode := "00001111";
						elsif Step = 1 then						-- Clock 1 till 2
							--DataI <= ReadResponse(1);
							RamDataToWrite := Operator(signed(ReadResponse(1)), signed(DataII), Operation);
							RamAddress := DestinationAddress;
							mode := "11110000";
							Step <= -1;
							Finish <= '1';
						end if;
							
					when Array_Alu =>
						DataII <= InPack(2);
						ArrayLength <= to_integer(unsigned(InPack(3)));
						DestinationAddress <= InPack(4);
						if to_integer(unsigned(InPack(3))) > 32 then
							Error <= '1';
						end if;
						
						if (Step > ArrayLength and Finish = '0')  then			-- Clock * size -> max 32
							mode := "11110000";
							RamDataToWrite := Operator(signed(ReadArray(ArrayIndPusher)), signed(DataII), Operation); -- Initail ArrayIndPusher = 0	
							RamAddress := byte((unsigned(DestinationAddress) + to_unsigned(ArrayIndPusher, 8)) mod 32);
							ArrayIndPusher <= ArrayIndPusher + 1;
							if ArrayIndPusher = (ArrayLength - 1) then
								Step <= -1;							-- Will + 1
								Finish <= '1';
								ArrayIndPusher <= 0;
							end if;
						else 
							if Step = 0 then							-- Clock * size -> max 32				
								--AddressI := InPack(1);
								ReadArray <= (others => (others => '0'));
								mode := "00001111";
							end if;
							if Step > 0 then 
								ReadArray(Step - 1) <= ReadResponse(1);
							end if;	
							RamAddress := byte((unsigned(InPack(1)) + to_unsigned(ArrayIndPusher, 8)) mod 32);
							ArrayIndPusher <= ArrayIndPusher + 1;
							if Step = ArrayLength then
								ArrayIndPusher <= 0;
							end if;
						end if;
						
					when Indirect_Addressing =>
						if Step = 0 then										-- Clock 0 till 1		
							DestinationAddress <= InPack(3);
							AddressI := InPack(1);
							RamAddress := AddressI;
							mode := "00001111";
						elsif Step = 1 then									-- Clock 1 till 2
							AddAddressII := InPack(2);
							DataI <= ReadResponse(1);
							mode := "00001111";
							RamAddress := AddAddressII;
						elsif Step = 2 then									-- Clock 2 till 3
							AddressII := ReadResponse(1);
							RamAddress := AddressII;
							mode := "00001111";	
						elsif Step = 3 then									-- Clock 3 till 4
							--DataII <= ReadResponse(1);
							RamDataToWrite := Operator(signed(DataI), signed(ReadResponse(1)), Operation);
							RamAddress := DestinationAddress;
							mode := "11110000";
							Step <= -1;										   -- Will + 1
							Finish <= '1';
						end if;
					when others =>
						Error <= '1';
				end case;
				Step <= Step + 1;
				SendToRam(0) <= mode;
				SendToRam(1) <= RamAddress;
				SendToRam(2) <= RamDataToWrite;
				SendToRam(3) <= (others => '0');
				SendToRam(4) <= (others => '0');
				SendToRam(5) <= (others => '0');
				SendToRam(6) <= (others => '0');
			end if;
		end if;
	end process;
	
end Behavioral;

